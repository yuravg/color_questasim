class class_a;
	int a
	function new();
	endfunction
endclass
